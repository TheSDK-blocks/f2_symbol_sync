../chisel/verilog/f2_symbol_sync.v